`timescale 1ns / 1ps

// -----------------------------------------------------------------------------
// Five-stage MIPS-like processor with automatic NOP insertion for load-use hazard
// -----------------------------------------------------------------------------
module proc (clk1, clk2);
input clk1, clk2;
// ------------------------ Pipeline Registers -------------------------------
reg [31:0] PC, IF_ID_IR, IF_ID_NPC;
reg [31:0] ID_EX_IR, ID_EX_NPC, ID_EX_A, ID_EX_B, ID_EX_Imm;
reg [2:0]  ID_EX_type, EX_MEM_type, MEM_WB_type;
reg [31:0] EX_MEM_IR, EX_MEM_ALUOut, EX_MEM_B;
reg        EX_MEM_cond;
reg [31:0] MEM_WB_IR, MEM_WB_ALUOut, MEM_WB_LMD;
// ----------------------------- Memories ------------------------------------
reg [31:0] Reg [0:31];
reg [31:0] Mem [0:1023];
// ----------------------------- Opcodes -------------------------------------
parameter ADD = 6'b000000, SUB = 6'b000001, AND = 6'b000010, OR  = 6'b000011,
          SLT = 6'b000100, MUL = 6'b000101, HLT = 6'b111111, LW  = 6'b001000,
          SW  = 6'b001001, ADDI= 6'b001010, SUBI= 6'b001011, SLTI= 6'b001100,
          BNEQZ=6'b001101, BEQZ=6'b001110,BEQ=6'b111110;
// --------------------------- Instruction Types -----------------------------
parameter RR_ALU = 3'b000, RM_ALU = 3'b001, LOAD = 3'b010, STORE = 3'b011,
          BRANCH = 3'b100, HALT  = 3'b101, NOP   = 3'b110;   // <- NEW
// ---------------------------- Flags ----------------------------------------
reg HALTED;
reg TAKEN_BRANCH;
reg STALL;                                           // <- NEW (load-use stall)

// ------------------------------ IF Stage -----------------------------------
always @ (posedge clk1) if (HALTED == 0) begin
     if (((EX_MEM_IR[31:26] == BEQZ) && (EX_MEM_cond == 1)) ||
                 ((EX_MEM_IR[31:26] == BNEQZ) && (EX_MEM_cond == 1))|| ((EX_MEM_IR[31:26] == BEQ) && (EX_MEM_cond == 1))) begin
        IF_ID_IR     <= Mem[EX_MEM_ALUOut];
        IF_ID_NPC    <= EX_MEM_ALUOut + 1;
        PC           <= EX_MEM_ALUOut + 1;
        TAKEN_BRANCH <= 1'b1;
    end else begin
        IF_ID_IR     <= Mem[PC];
        IF_ID_NPC    <= PC + 1;
        PC           <= PC + 1;
    end
end

// ------------------------------ ID Stage -----------------------------------
always @ (posedge clk2) if (HALTED == 0) begin
        // Normal decode operations
        ID_EX_NPC  <= IF_ID_NPC;
        ID_EX_IR   <= IF_ID_IR;
        ID_EX_Imm  <= {{16{IF_ID_IR[15]}}, IF_ID_IR[15:0]};
        // -------------------- Register Read / Forwarding ------------------
        // Forward A
        if (( EX_MEM_type == RM_ALU ) && // rm 1st operand
            (EX_MEM_IR[20:16] == IF_ID_IR[25:21]) && (IF_ID_IR[25:21] != 0))
            begin
            ID_EX_A <=  EX_MEM_ALUOut;
            end
            else if(( EX_MEM_type == RR_ALU ) &&
            (EX_MEM_IR[15:11] == IF_ID_IR[25:21]) && (IF_ID_IR[25:21] != 0))
            begin
            ID_EX_A <=  EX_MEM_ALUOut;
            end
           else if (( EX_MEM_type == LOAD ) &&
            (EX_MEM_IR[20:16] == IF_ID_IR[25:21]) && (IF_ID_IR[25:21] != 0))
            begin
            ID_EX_A <=  Mem[EX_MEM_ALUOut] ;
            end
        else
        begin
            ID_EX_A <= (IF_ID_IR[25:21] == 0) ? 0 : Reg[IF_ID_IR[25:21]];
            end
        // Forward B
        if (( EX_MEM_type == RM_ALU ) &&
            (EX_MEM_IR[20:16] == IF_ID_IR[20:16]) && (IF_ID_IR[20:16] != 0))
            begin
            ID_EX_B <= (EX_MEM_type == LOAD) ?  Mem[EX_MEM_ALUOut] : EX_MEM_ALUOut;
            end
            else if(( EX_MEM_type == RR_ALU ) &&
            (EX_MEM_IR[15:11] == IF_ID_IR[20:16]) && (IF_ID_IR[20:16] != 0))
            begin
            ID_EX_B <= (EX_MEM_type == LOAD) ?  Mem[EX_MEM_ALUOut] : EX_MEM_ALUOut;
            end
            else if (( EX_MEM_type == LOAD ) &&
            (EX_MEM_IR[20:16] == IF_ID_IR[20:16]) && (IF_ID_IR[20:16] != 0))
            begin
            ID_EX_B <= (EX_MEM_type == LOAD) ?  Mem[EX_MEM_ALUOut] : EX_MEM_ALUOut;
            end
        else
        begin
            ID_EX_B <= (IF_ID_IR[20:16] == 0) ? 0 : Reg[IF_ID_IR[20:16]];
            end
        // Instruction type
        case (IF_ID_IR[31:26])
            ADD, SUB, AND, OR, SLT, MUL: ID_EX_type <= RR_ALU;
            ADDI, SUBI, SLTI:            ID_EX_type <= RM_ALU;
            LW:                          ID_EX_type <= LOAD;
            SW:                          ID_EX_type <= STORE;
            BNEQZ,BEQZ ,BEQ:              ID_EX_type <= BRANCH;
            HLT:                         ID_EX_type <= HALT;
            default:                     ID_EX_type <= NOP;
        endcase
    end

// ------------------------------ EX Stage -----------------------------------
always @ (posedge clk1) if (HALTED == 0) begin
    EX_MEM_type <= ID_EX_type;
    EX_MEM_IR   <= ID_EX_IR;
    TAKEN_BRANCH <= 0;
    case (ID_EX_type)
        NOP: EX_MEM_ALUOut <= 0;
        RR_ALU: begin
            case (ID_EX_IR[31:26])
                ADD: EX_MEM_ALUOut <= ID_EX_A + ID_EX_B;
                SUB: EX_MEM_ALUOut <= ID_EX_A - ID_EX_B;
                AND: EX_MEM_ALUOut <= ID_EX_A & ID_EX_B;
                OR:  EX_MEM_ALUOut <= ID_EX_A | ID_EX_B;
                SLT: EX_MEM_ALUOut <= (ID_EX_A < ID_EX_B);
                MUL: EX_MEM_ALUOut <= ID_EX_A * ID_EX_B;
                default: EX_MEM_ALUOut <= 32'hxxxx_xxxx;
            endcase
        end
        RM_ALU: begin
            case (ID_EX_IR[31:26])
                ADDI: EX_MEM_ALUOut <= ID_EX_A + ID_EX_Imm;
                SUBI: EX_MEM_ALUOut <= ID_EX_A - ID_EX_Imm;
                SLTI: EX_MEM_ALUOut <= (ID_EX_A < ID_EX_Imm);
                default: EX_MEM_ALUOut <= 32'hxxxx_xxxx;
            endcase
        end
        LOAD, STORE: begin
            EX_MEM_ALUOut <= ID_EX_A + ID_EX_Imm;
            EX_MEM_B      <= ID_EX_B;
        end
        BRANCH: begin
            case (ID_EX_IR[31:26])
                BEQZ: begin 
                    EX_MEM_ALUOut <= ID_EX_NPC + ID_EX_Imm;
                    EX_MEM_cond   <= (ID_EX_A == 0);
                end
                BNEQZ: begin 
                    EX_MEM_ALUOut <= ID_EX_NPC + ID_EX_Imm;
                    EX_MEM_cond   <= (ID_EX_A != 0);
                end
                BEQ: begin 
                    EX_MEM_ALUOut <= ID_EX_NPC + ID_EX_Imm;
                    EX_MEM_cond   <= (ID_EX_A == ID_EX_B);
                end
                default: begin
                    EX_MEM_ALUOut <= 32'hxxxx_xxxx;
                    EX_MEM_cond <= 1'bx;
                end
            endcase
        end
    endcase
end


// ------------------------------ MEM Stage ----------------------------------
always @ (posedge clk2) 
    if (HALTED == 0) begin
        MEM_WB_type <= EX_MEM_type;
        MEM_WB_IR   <= EX_MEM_IR;

        case (EX_MEM_type)
            RR_ALU, RM_ALU: MEM_WB_ALUOut <= EX_MEM_ALUOut;
            LOAD:           MEM_WB_LMD    <= Mem[EX_MEM_ALUOut];
            STORE:          if (TAKEN_BRANCH == 0)
                                Mem[EX_MEM_ALUOut] <= EX_MEM_B;
            // NOP and others do nothing
        endcase
    end


// ------------------------------ WB Stage -----------------------------------
always @ (posedge clk1) 
begin
    if (TAKEN_BRANCH == 0) begin
        case (MEM_WB_type)
            RR_ALU: Reg[MEM_WB_IR[15:11]] <= MEM_WB_ALUOut;
            RM_ALU: Reg[MEM_WB_IR[20:16]] <= MEM_WB_ALUOut;
            LOAD:   Reg[MEM_WB_IR[20:16]] <= MEM_WB_LMD;
            HALT:   HALTED <= 1'b1;
            default: ; // NOP has no effect
        endcase
    end
end

endmodule